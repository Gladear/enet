module enet

fn C.enet_initialize() int

fn C.enet_deinitialize()
