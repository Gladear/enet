module enet

pub type Compressor = C._ENetCompressor
